`ifndef PARAMS_H_
`define PARAMS_H_

`define n_BIT_CLKS_9600    2500 // 24MHz / 9600baud
`define n_BIT_CLKS_230400  104  // 24MHz / 230400baud

`define n_BIT_CLKS `n_BIT_CLKS_230400

`endif